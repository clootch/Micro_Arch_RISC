module memory(
	
);
endmodule