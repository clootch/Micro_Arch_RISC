module memory(
	
);